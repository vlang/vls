import vls

const = (
	sample = '
module main

fn main() {
	println(\'foo\')
}
	'
)

fn test_position_to_lsp_pos() {
	// TODO:
}

fn test_position_to_lsp_range() {
	// TODO:
}

fn test_compute_offset() {
	// TODO:
}