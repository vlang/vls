module log

fn test_notification_send() {
	
}