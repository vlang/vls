module vls

const (
	v_exec_name   = 'v.exe'
	path_list_sep = ';'
)
