module def

pub fn hello() {}