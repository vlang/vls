module abc

pub struct Def {}