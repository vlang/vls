module abc

pub struct Point {
	a int
	b int
}

pub fn this_is_a_function() string {
	return 'wee'
}