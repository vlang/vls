// TODO: This code will be probably moved to features.v depending on the
// complexity of the code. What you're seeing here is not final so please
// bear in mind about it. 
// TODO: Add tests for it
module vls

import lsp
import os
import jsonrpc
import json
import v.ast
import v.table

struct CompletionItemConfig {
mut:
	pub_only            bool = true
	file                ast.File
	offset              int
	table               &table.Table
	show_global         bool = true
	show_only_global_fn bool
	show_local          bool       = true
	filter_type         table.Type = table.Type(0)
	fields_only         bool
	file_imports        []string
}

fn (mut cfg CompletionItemConfig) completion_items_from_stmt(stmt ast.Stmt) []lsp.CompletionItem {
	mut completion_items := []lsp.CompletionItem{}
	match stmt {
		ast.ExprStmt {
			completion_items << cfg.completion_items_from_expr(stmt.expr)
		}
		ast.AssignStmt {
			if stmt.op != .decl_assign {
				cfg.show_global = false
				cfg.show_only_global_fn = false
				cfg.filter_type = stmt.left_types[stmt.left_types.len - 1]
			}
		}
		ast.Import {
			dir := os.dir(cfg.file.path)
			dir_contents := os.ls(dir) or { []string{} }
			// list all folders
			completion_items << cfg.completion_items_from_dir(dir, dir_contents)
			// list all vlib
			// TODO: vlib must be computed at once only
		}
		else {}
	}
	return completion_items
}

fn (mut cfg CompletionItemConfig) completion_items_from_table(prefix_name string) []lsp.CompletionItem {
	mut completion_items := []lsp.CompletionItem{}
	if cfg.show_global && cfg.show_only_global_fn {
		return completion_items
	}
	for sym_name, idx in cfg.table.type_idxs {
		if idx <= 0 || idx >= cfg.table.types.len || !sym_name.starts_with('${prefix_name}.') {
			continue
		}
		type_sym := unsafe { &cfg.table.types[idx] }
		completion_items <<
			cfg.completion_items_from_type_info(sym_name.all_after('${prefix_name}.'), type_sym.info, false)
	}
	return completion_items
}

fn (mut cfg CompletionItemConfig) completion_items_from_expr(expr ast.Expr) []lsp.CompletionItem {
	mut completion_items := []lsp.CompletionItem{}
	mut expr_type := table.Type(0)
	// TODO: support for infix/postfix expr
	match expr {
		ast.SelectorExpr {
			expr_type = expr.expr_type
			if expr_type == 0 && expr.expr is ast.Ident {
				ident := expr.expr as ast.Ident
				if ident.name !in cfg.file_imports {
					return completion_items
				}
				// NB: symbols of the said module does not show the full list
				// unless by pressing cmd/ctrl+space or by pressing escape key
				// + deleting the dot + typing again the dot
				completion_items << cfg.completion_items_from_table(ident.name)
				for _, fnn in cfg.table.fns {
					if fnn.mod != ident.name || !fnn.is_pub {
						continue
					}
					completion_items << cfg.completion_items_from_fn(fnn, false)
				}
			} else if expr_type != 0 {
				type_sym := cfg.table.get_type_symbol(expr_type)
				completion_items <<
					cfg.completion_items_from_type_info('', type_sym.info, true)
				if type_sym.kind == .array || type_sym.kind == .map {
					base_symbol_name := if type_sym.kind == .array { 'array' } else { 'map' }
					if base_type_sym := cfg.table.find_type(base_symbol_name) {
						completion_items <<
							cfg.completion_items_from_type_info('', base_type_sym.info, true)
					}
				}
				// list all methods
				for m in type_sym.methods {
					completion_items << cfg.completion_items_from_fn(m, true)
				}
			}
			return completion_items
		}
		ast.CallExpr {
			current_arg_idx := expr.args.len
			if current_arg_idx < expr.expected_arg_types.len {
				cfg.show_local = true
				cfg.show_global = false
				cfg.filter_type = expr.expected_arg_types[current_arg_idx]
			} else {
				cfg.show_local = false
				cfg.show_global = false
			}
			return completion_items
		}
		ast.StructInit {
			cfg.show_global = false
			cfg.show_local = false
			field_node := find_ast_by_pos(expr.fields.map(ast.Node(it)), cfg.offset - 1) or {
				ast.Node{}
			}
			if field_node is ast.StructInitField {
				// NB: enable local results only if the node is a field
				cfg.show_local = true
				field_type_sym := cfg.table.get_type_symbol(field_node.expected_type)
				completion_items <<
					cfg.completion_items_from_type_info('', field_type_sym.info, field_type_sym.info is table.Enum)
				cfg.filter_type = field_node.expected_type
			} else {
				// if structinit is empty or not within the field position, 
				// it must show the list of missing fields instead
				defined_fields := expr.fields.map(it.name)
				struct_type_sym := cfg.table.get_type_symbol(expr.typ)
				struct_type_info := struct_type_sym.info as table.Struct
				for field in struct_type_info.fields {
					if field.name in defined_fields {
						continue
					}
					completion_items << lsp.CompletionItem{
						label: '$field.name:'
						kind: .field
						insert_text: '$field.name: \$0'
						insert_text_format: .snippet
					}
				}
			}
		}
		else {}
	}
	return completion_items
}

fn (mut cfg CompletionItemConfig) completion_items_from_fn(fnn table.Fn, is_method bool) lsp.CompletionItem {
	mut i := 0
	mut insert_text := fnn.name.all_after(fnn.mod + '.')
	kind := if is_method { lsp.CompletionItemKind.method } else { lsp.CompletionItemKind.function }
	if fnn.is_generic {
		insert_text += '<\${$i:T}>'
	}
	insert_text += '('
	for j, param in fnn.params {
		if is_method && j == 0 {
			continue
		}
		i++
		insert_text += '\${$i:$param.name}'
		if j < fnn.params.len - 1 {
			insert_text += ', '
		}
	}
	insert_text += ')'
	if fnn.return_type.has_flag(.optional) {
		insert_text += ' or { panic(err) }'
	}
	return lsp.CompletionItem{
		label: fnn.name.all_after(fnn.mod + '.')
		kind: kind
		insert_text_format: .snippet
		insert_text: insert_text
	}
}

fn (mut cfg CompletionItemConfig) completion_items_from_type_info(name string, type_info table.TypeInfo, fields_only bool) []lsp.CompletionItem {
	mut completion_items := []lsp.CompletionItem{}
	match type_info {
		table.Struct {
			if !fields_only {
				mut insert_text := '$name{\n'
				mut i := type_info.fields.len - 1
				for field in type_info.fields {
					if field.has_default_expr {
						continue
					}
					insert_text += '\t$field.name: \$$i\n'
					i--
				}
				insert_text += '}'
				completion_items << lsp.CompletionItem{
					label: '$name{}'
					kind: .struct_
					insert_text: insert_text
					insert_text_format: .snippet
				}
			} else {
				for field in type_info.fields {
					completion_items << lsp.CompletionItem{
						label: field.name
						kind: .field
						insert_text: field.name
					}
				}
			}
		}
		table.Enum {
			for val in type_info.vals {
				label := if fields_only { '.$val' } else { '${name}.$val' }
				completion_items << lsp.CompletionItem{
					label: label
					kind: .enum_member
					insert_text: label
				}
			}
		}
		table.Alias, table.SumType, table.FnType, table.Interface {
			completion_items << lsp.CompletionItem{
				label: name
				kind: .type_parameter
				insert_text: name
			}
		}
		else {}
	}
	return completion_items
}

fn (cfg CompletionItemConfig) completion_items_from_dir(dir string, dir_contents []string) []lsp.CompletionItem {
	mut completion_items := []lsp.CompletionItem{}
	for name in dir_contents {
		full_path := os.join_path(dir, name)
		if !os.is_dir(full_path) || name in cfg.file_imports {
			continue
		}
		subdir_contents := os.ls(full_path) or { []string{} }
		completion_items << cfg.completion_items_from_dir(full_path, subdir_contents)
		if name == 'modules' {
			continue
		}
		completion_items << lsp.CompletionItem{
			label: name
			kind: .folder
			insert_text: name
		}
	}
	return completion_items
}

// TODO: make params use lsp.CompletionParams in the future
fn (mut ls Vls) completion(id int, params string) {
	completion_params := json.decode(lsp.CompletionParams, params) or { panic(err) }
	file_uri := completion_params.text_document.uri
	file := ls.files[file_uri.str()]
	src := ls.sources[file_uri.str()]
	mut pos := completion_params.position
	mut ctx := completion_params.context
	mut completion_items := []lsp.CompletionItem{}
	mut cfg := CompletionItemConfig{
		file: file
		file_imports: file.imports.map(if it.alias.len > 0 { it.alias } else { it.mod })
		offset: compute_offset(src, pos.line, pos.character)
		table: ls.tables[os.dir(file_uri)]
	}
	// adjust context data if the trigger symbols are on the left
	if ctx.trigger_kind == .invoked && cfg.offset - 1 >= 0 && file.stmts.len > 0 && src.len > 3 {
		if src[cfg.offset - 1] in [`.`, `:`, `=`, `{`, `,`, `(`] {
			ctx = lsp.CompletionContext{
				trigger_kind: .trigger_character
				trigger_character: src[cfg.offset - 1].str()
			}
		} else if src[cfg.offset - 1] == ` ` &&
			cfg.offset - 2 >= 0 && src[cfg.offset - 2] !in [src[cfg.offset - 1], `.`] {
			ctx = lsp.CompletionContext{
				trigger_kind: .trigger_character
				trigger_character: src[cfg.offset - 2].str()
			}
			cfg.offset -= 2
			pos = {
				pos |
				character: pos.character - 2
			}
		}
	}
	if ctx.trigger_kind == .trigger_character {
		if ctx.trigger_character == '.' && (cfg.offset - 1 >= 0 && src[cfg.offset - 1] != ` `) {
			cfg.show_global = false
			cfg.show_local = false
			cfg.offset -= 2
		}
		node := find_ast_by_pos(file.stmts.map(ast.Node(it)), cfg.offset) or { ast.Node{} }
		if node is ast.Stmt {
			completion_items << cfg.completion_items_from_stmt(node)
		} else if node is ast.Expr {
			completion_items << cfg.completion_items_from_expr(node)
		}
	} else if ctx.trigger_kind == .invoked && (file.stmts.len == 0 || src.len <= 3) {
		// should never happen but just to make sure
		cfg.show_global = false
		cfg.show_local = false
		folder_name := os.base(os.dir(file_uri.str())).replace(' ', '_')
		module_name_suggestions := ['module main', 'module $folder_name']
		for sg in module_name_suggestions {
			completion_items << lsp.CompletionItem{
				label: sg
				insert_text: sg
				kind: .variable
			}
		}
	} else {
		cfg.show_only_global_fn = true
	}
	if cfg.show_local {
		if cfg.filter_type == 0 {
			// get the module names
			for imp in file.imports {
				if imp.mod in ls.invalid_imports[file_uri.str()] {
					continue
				}
				completion_items << lsp.CompletionItem{
					label: if imp.alias.len > 0 {
						imp.alias
					} else {
						imp.mod
					}
					kind: .module_
				}
			}
		}
		inner_scope := file.scope.innermost(cfg.offset)
		for scope in [file.scope, inner_scope] {
			for _, obj in scope.objects {
				mut name := ''
				match obj {
					ast.ConstField, ast.Var {
						if cfg.filter_type != 0 && obj.typ != cfg.filter_type {
							continue
						}
						name = obj.name
					}
					else {
						continue
					}
				}
				mut kind := lsp.CompletionItemKind.variable
				if obj is ast.ConstField {
					name = name.all_after('${obj.mod}.')
					kind = .constant
				}
				completion_items << lsp.CompletionItem{
					label: name
					kind: kind
					insert_text: name
				}
			}
		}
	}
	if cfg.show_global {
		completion_items << cfg.completion_items_from_table(file.mod.name)
		// include functions from builtin and within the same namespace
		for _, fnn in cfg.table.fns {
			if (fnn.mod == 'builtin' &&
				fnn.name in ls.builtin_symbols) ||
				(fnn.mod == file.mod.name && fnn.name != 'main.main') {
				completion_items << cfg.completion_items_from_fn(fnn, false)
			}
		}
	}
	ls.send(json.encode(jsonrpc.Response<[]lsp.CompletionItem>{
		id: id
		result: completion_items
	}))
	unsafe { completion_items.free() }
}
