module main

fn test_compilation() {
	println('ok')
	assert true
}
