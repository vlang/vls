module lsp

// method: ‘textDocument/definition’
// response: Location | []Location | []LocationLink | none
// request: TextDocumentPositionParams

// method: ‘textDocument/typeDefinition’
// response: Location | []Location | []LocationLink | none
// request: TextDocumentPositionParams