module vls

const (
	v_exec_name = 'v'
	path_list_sep = ':'
)
