module abc