module ghi

pub fn world() {}