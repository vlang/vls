module vls


fn (ls Vls) did_change_watched_files(id int, params string) string {

}
