module errors

pub const (
	unknown_node_type_error               = 'unknown_node_type_error'
	bool_string_cast_error                = 'bool_string_cast_error'
	constant_mutation_error               = 'constant_mutation_error'
	decomposition_error                   = 'decomposition_error'
	defer_break_error                     = 'defer_break_error'
	empty_enum_error                      = 'empty_enum_error'
	enum_default_value_error              = 'enum_default_value_error'
	enum_duplicate_member_error           = 'enum_duplicate_member_error'
	enum_duplicate_value_error            = 'enum_duplicate_value_error'
	enum_value_overflow_error             = 'enum_value_overflow_error'
	unexpected_argument_error_single      = 'unexpected_argument_error_single'
	unexpected_argument_error_plural      = 'unexpected_argument_error_plural'
	float_modulo_error                    = 'float_modulo_error'
	match_duplicate_branch_error          = 'match_duplicate_branch_error'
	match_invalid_case_value_error        = 'match_invalid_case_value_error'
	match_invalid_sumtype_variant_error   = 'match_invalid_sumtype_variant_error'
	match_expr_no_expression_value_error  = 'match_expr_no_expression_value_error'
	match_expr_value_type_mismatch        = 'match_expr_value_type_mismatch'
	match_range_value_type_mismatch       = 'match_range_value_type_mismatch'
	match_sumtype_not_exhaustive_error    = 'match_sumtype_not_exhaustive_error'
	mismatched_type_error                 = 'mismatched_type_error'
	nonloop_break_error                   = 'nonloop_break_error'
	not_found_error                       = 'not_found_error'
	not_public_error                      = 'not_public_error'
	non_reference_return_error            = 'non_reference_return_error'
	if_expr_non_bool_cond_error           = 'if_expr_non_bool_cond_error'
	if_expr_no_else_error                 = 'if_expr_no_else_error'
	if_no_expression_value_error          = 'if_no_expression_value_error'
	imaginary_mutation_error              = 'imaginary_mutation_error'
	immutable_variable_error              = 'immutable_variable_error'
	invalid_argument_error                = 'invalid_argument_error'
	invalid_option_propagate_call_error   = 'invalid_option_propagate_call_error'
	undefined_ident_assignment_error      = 'undefined_ident_assignment_error'
	undefined_operation_error             = 'undefined_operation_error'
	unhandled_optional_fn_call_error      = 'unhandled_optional_fn_call_error'
	unhandled_optional_selector_error     = 'unhandled_optional_selector_error'
	unknown_type_error                    = 'unknown_type_error'
	unknown_function_error                = 'unknown_function_error'
	unknown_field_error                   = 'unknown_field_error'
	unknown_method_or_field_error         = 'unknown_method_or_field_error'
	uninitialized_reference_field_error   = 'uninitialized_reference_field_error'
	ambiguous_method_error                = 'ambiguous_method_error'
	ambiguous_field_error                 = 'ambiguous_field_error'
	ambiguous_call_error                  = 'ambiguous_call_error'
	append_type_mismatch_error            = 'append_type_mismatch_error'
	array_append_expr_error               = 'array_append_expr_error'
	invalid_array_element_type_error      = 'invalid_array_element_type_error'
	invalid_enum_casting_error            = 'invalid_enum_casting_error'
	invalid_sumtype_array_init_error      = 'invalid_sumtype_array_init_error'
	invalid_assignment_error              = 'invalid_assignment_error'
	invalid_return_error                  = 'invalid_return_error'
	selective_const_import_error          = 'selective_const_import_error'
	send_channel_invalid_chan_type_error  = 'send_channel_invalid_chan_type_error'
	send_channel_invalid_value_type_error = 'send_channel_invalid_value_type_error'
	send_operator_in_var_decl_error       = 'send_operator_in_var_decl_error'
	invalid_assert_type_error             = 'invalid_assert_type_error'
	invalid_void_return_error             = 'invalid_void_return_error'
	typedef_map_init_error                = 'typedef_map_init_error'
	unnecessary_if_parenthesis_error      = 'unnecessary_if_parenthesis_error'
	unreachable_code_error                = 'unreachable_code_error'
	untyped_empty_array_error             = 'untyped_empty_array_error'
	unused_expression_error               = 'unused_identifier_error'
	unwrapped_option_binary_expr_error    = 'unwrapped_option_binary_expr_error'
	unexpected_return_error               = 'unexpected_return_error'
	void_value_return_error               = 'void_value_return_error'
	void_symbol_casting_error             = 'void_symbol_casting_error'
	wrong_error_propagation_error         = 'wrong_error_propagation_error'
)

pub const message_templates = {
	unknown_node_type_error:               'unknown node `%s`'
	bool_string_cast_error:                'cannot cast type `bool` to string, use `%s.str()` instead.'
	constant_mutation_error:               'cannot modify constant `%s`'
	decomposition_error:                   'decomposition can only be used on arrays'
	defer_break_error:                     '`break` is not allowed in defer statements'
	empty_enum_error:                      'enum cannot be empty'
	enum_default_value_error:              'default value for enum has to be an integer'
	enum_duplicate_member_error:           'field name `%s` duplicate'
	enum_duplicate_value_error:            'enum value `%s` already exists'
	enum_value_overflow_error:             'enum value overflows'
	unexpected_argument_error_plural:      'expected %s arguments, but got %s'
	unexpected_argument_error_single:      'expected %s argument, but got %s'
	float_modulo_error:                    'float modulo not allowed, use math.fmod() instead'
	match_duplicate_branch_error:          'match case `%s` is handled more than once'
	match_invalid_case_value_error:        'cannot match `%s` with `%s`'
	match_invalid_sumtype_variant_error:   '`%` has no variant `%s`'
	match_expr_no_expression_value_error:  '`match` expression requires an expression as the last statement of every branch'
	match_expr_value_type_mismatch:        'return type mismatch, it should be `%s`'
	match_range_value_type_mismatch:       'mismatched range types'
	match_sumtype_not_exhaustive_error:    r'match must be exhaustive (add match branches for {types} or `else {}` at the end)'
	mismatched_type_error:                 'mismatched types `%s` and `%s`'
	nonloop_break_error:                   'break statement not within a loop'
	not_found_error:                       'symbol `%s` not found'
	not_public_error:                      'symbol `%s` not public'
	non_reference_return_error:            'fn `%s` expects you to return a reference type `%s`, but you are returning `%s` instead'
	if_expr_non_bool_cond_error:           'non-bool type `%s` used as if condition'
	if_expr_no_else_error:                 '`if` expression needs `else` clause'
	if_no_expression_value_error:          '`if` expression requires an expression as the last statement of every branch'
	imaginary_mutation_error:              'cannot modify blank `_` identifier'
	immutable_variable_error:              '`%s` is immutable, declare it with `mut` to make it mutable'
	invalid_argument_error:                'cannot use `%s` as `%s` in argument %s to `%s`'
	invalid_option_propagate_call_error:   'unexpected `?`, the function `%s` does neither return an optional nor a result'
	undefined_ident_assignment_error:      'undefined ident: `%s` (use `:=` to declare a variable)'
	undefined_operation_error:             'undefined operation `%s` %s `%s`'
	unhandled_optional_fn_call_error:      '%s() returns an option, so it should have either an `or {}` block, or `?` at the end'
	unhandled_optional_selector_error:     'cannot access fields of an optional, handle the error with `or {...}` or propagate it with `?`'
	unknown_type_error:                    'unknown type `%s`'
	unknown_function_error:                'unknown function: %s'
	unknown_field_error:                   'type `%s` has no field named `%s`'
	unknown_method_or_field_error:         'unknown method or field: `%s.%s`'
	uninitialized_reference_field_error:   'reference field `%s.%s` must be initialized'
	ambiguous_method_error:                'ambiguous method `%s`'
	ambiguous_field_error:                 'ambiguous field `%s`'
	ambiguous_call_error:                  'ambiguous call to: `%s`, may refer to fn `%s` or variable `%s`'
	append_type_mismatch_error:            'cannot append `%s` to `%s`'
	array_append_expr_error:               'array append cannot be used in an expression'
	invalid_array_element_type_error:      'invalid array element: expected `%s`, not `%s`'
	invalid_enum_casting_error:            '%s does not represent a value of enum %s'
	invalid_sumtype_array_init_error:      'cannot initialize sum type array without default value'
	invalid_return_error:                  'cannot use `%s` as type `%s` in return argument'
	invalid_void_return_error:             'expected `%s` argument'
	send_channel_invalid_chan_type_error:  'cannot push on non-channel `%s`'
	invalid_assignment_error:              'cannot assign to `%s`: expected `%s`, not `%s`'
	selective_const_import_error:          r'cannot selective import constant `{{var}}` from `{{module}}`, import `{{module}}` and use `{{module}}.{{var}}` instead'
	send_channel_invalid_value_type_error: 'cannot push `%s` on `%s`'
	send_operator_in_var_decl_error:       '<- operator can only be used with `chan` types'
	invalid_assert_type_error:             'assert can be used only with `bool` expressions, but found `%s` instead'
	typedef_map_init_error:                r'direct map alias init is not possible, use `{{type_name}}({{map_type}}{})` instead'
	unnecessary_if_parenthesis_error:      'unnecessary `()` in `if` condition, use `if expr {` instead of `if (expr) {`'
	unreachable_code_error:                'unreachable code'
	untyped_empty_array_error:             'array_init: no type specified (maybe: `[]Type{}` instead of `[]`)'
	unused_expression_error:               '`%s` evaluated but not used'
	unwrapped_option_binary_expr_error:    'unwrapped optional cannot be used in an infix expression'
	unexpected_return_error:               'unexpected argument, current function does not return anything'
	void_value_return_error:               '`%s` used as value'
	void_symbol_casting_error:             'expression does not return a value so it cannot be cast'
	wrong_error_propagation_error:         'to propagate the optional call, `%s` must return an optional'
}
