module def

pub fn hello() string {
	return 'hello'
}