module efg

pub struct Vector {
	x int
	y int
}