module gfx

[typedef]
pub struct C.Foo {
	bar   int
	baz   string
	data  voidptr
	count int
}
